library verilog;
use verilog.vl_types.all;
entity extensor_sinal_vlg_vec_tst is
end extensor_sinal_vlg_vec_tst;
