LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY mux4to1_64 IS PORT(
	IN0,IN1,IN2,IN3: IN STD_LOGIC_VECTOR (63 DOWNTO 0);
	SEL : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
	S : OUT STD_LOGIC_VECTOR (63 DOWNTO 0)
);
END ENTITY;
	
ARCHITECTURE projeto OF mux4to1_64 IS
BEGIN
S <=	IN3 WHEN SEL = "11" ELSE
		IN2 WHEN SEL = "10" ELSE
		IN1 WHEN SEL = "01" ELSE
		IN0;
END projeto;
