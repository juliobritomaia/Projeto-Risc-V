LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY mux2to1_64 IS PORT(
	IN0,IN1 : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
	SEL : IN STD_LOGIC;
	S : OUT STD_LOGIC_VECTOR (63 DOWNTO 0)
);
END ENTITY;
	
ARCHITECTURE projeto OF mux2to1_64 IS
BEGIN
S <=	IN1 WHEN SEL = '1' ELSE
		IN0;
END projeto;
